library work;
  use work.globals.all;

package zeta_lut is

  type zeta_array_t is array (0 to n - 1) of modq_t;

  -- constant zetas : zeta_array_t :=
  -- (
  --   0 => 1,
  --   1 => 42,
  --   2 => 69,
  --   3 => 73,
  --   4 => 15,
  --   5 => 65,
  --   6 => 18,
  --   7 => 78
  -- );

  constant zetas : zeta_array_t :=
  (
    0   => 4193792,
    1   => 2091667,
    2   => 4450022,
    3   => 7100756,
    4   => 2706023,
    5   => 342297,
    6   => 5037034,
    7   => 5341501,
    8   => 2725464,
    9   => 900702,
    10  => 3412210,
    11  => 6366809,
    12  => 6681150,
    13  => 4613401,
    14  => 189548,
    15  => 5441381,
    16  => 1826347,
    17  => 266997,
    18  => 7122806,
    19  => 7838005,
    20  => 4519302,
    21  => 2842341,
    22  => 4656075,
    23  => 7953734,
    24  => 6262231,
    25  => 7725090,
    26  => 7709315,
    27  => 5196991,
    28  => 811944,
    29  => 7047359,
    30  => 1285669,
    31  => 7826001,
    32  => 237124,
    33  => 5037939,
    34  => 6927966,
    35  => 1500165,
    36  => 6718724,
    37  => 3437287,
    38  => 44288,
    39  => 2213111,
    40  => 7830929,
    41  => 495491,
    42  => 5412772,
    43  => 1957272,
    44  => 3507263,
    45  => 5386378,
    46  => 5971092,
    47  => 183443,
    48  => 3119733,
    49  => 4860065,
    50  => 5190273,
    51  => 5796124,
    52  => 3539968,
    53  => 4055324,
    54  => 2389356,
    55  => 6712985,
    56  => 1757237,
    57  => 4823422,
    58  => 7998430,
    59  => 810149,
    60  => 3900724,
    61  => 7929317,
    62  => 5361315,
    63  => 3937738,
    64  => 5771523,
    65  => 2316500,
    66  => 4702672,
    67  => 5834105,
    68  => 3077325,
    69  => 5942594,
    70  => 508951,
    71  => 3866901,
    72  => 7300517,
    73  => 909542,
    74  => 2147896,
    75  => 2454455,
    76  => 3505694,
    77  => 2635921,
    78  => 3159746,
    79  => 7959518,
    80  => 8021166,
    81  => 7144689,
    82  => 4296819,
    83  => 6709241,
    84  => 3574422,
    85  => 5790267,
    86  => 1653064,
    87  => 6577327,
    88  => 6980856,
    89  => 2031748,
    90  => 8357436,
    91  => 1616392,
    92  => 954230,
    93  => 5062207,
    94  => 7567685,
    95  => 8332111,
    96  => 7504169,
    97  => 5933984,
    98  => 2176455,
    99  => 2235880,
    100 => 5842901,
    101 => 1735879,
    102 => 904516,
    103 => 1717735,
    104 => 2619752,
    105 => 8337157,
    106 => 7969390,
    107 => 185531,
    108 => 6779997,
    109 => 1903435,
    110 => 1315589,
    111 => 1612842,
    112 => 3111497,
    113 => 7183191,
    114 => 4747489,
    115 => 594136,
    116 => 2348700,
    117 => 2486353,
    118 => 759969,
    119 => 8119771,
    120 => 4010497,
    121 => 7611795,
    122 => 1852771,
    123 => 4686184,
    124 => 2071892,
    125 => 3306115,
    126 => 4751448,
    127 => 7534263,
    128 => 25847,
    129 => 3407706,
    130 => 6851714,
    131 => 1917081,
    132 => 95776,
    133 => 286988,
    134 => 264944,
    135 => 3523897,
    136 => 1024112,
    137 => 1859098,
    138 => 7396998,
    139 => 2432395,
    140 => 6736599,
    141 => 1250494,
    142 => 4827145,
    143 => 6144432,
    144 => 2353451,
    145 => 2434439,
    146 => 1939314,
    147 => 5548557,
    148 => 5336701,
    149 => 2691481,
    150 => 8371839,
    151 => 1723600,
    152 => 4520680,
    153 => 5257975,
    154 => 7151892,
    155 => 162844,
    156 => 531354,
    157 => 1237275,
    158 => 6795489,
    159 => 3919660,
    160 => 7602457,
    161 => 2244091,
    162 => 3475950,
    163 => 777191,
    164 => 4788269,
    165 => 5038140,
    166 => 7280319,
    167 => 7404533,
    168 => 7260833,
    169 => 6767243,
    170 => 4686924,
    171 => 3369112,
    172 => 6239768,
    173 => 1869119,
    174 => 8202977,
    175 => 7403526,
    176 => 5495562,
    177 => 4621053,
    178 => 5223087,
    179 => 4656147,
    180 => 8079950,
    181 => 1247620,
    182 => 8169440,
    183 => 7276084,
    184 => 8360995,
    185 => 7855319,
    186 => 1349076,
    187 => 1652634,
    188 => 5823537,
    189 => 1312455,
    190 => 4499357,
    191 => 1400424,
    192 => 7861508,
    193 => 3817976,
    194 => 5339162,
    195 => 7005614,
    196 => 3530437,
    197 => 4108315,
    198 => 3097992,
    199 => 269760,
    200 => 3585928,
    201 => 819034,
    202 => 2715295,
    203 => 8215696,
    204 => 4558682,
    205 => 4832145,
    206 => 6529015,
    207 => 6094090,
    208 => 6288512,
    209 => 3513181,
    210 => 7380215,
    211 => 6533464,
    212 => 5512770,
    213 => 1265009,
    214 => 5130689,
    215 => 1910376,
    216 => 5102745,
    217 => 3207046,
    218 => 7072248,
    219 => 3014001,
    220 => 3881043,
    221 => 6950192,
    222 => 6940675,
    223 => 7018208,
    224 => 466468,
    225 => 4817955,
    226 => 6795196,
    227 => 3406031,
    228 => 3915439,
    229 => 203044,
    230 => 3958618,
    231 => 472078,
    232 => 6271868,
    233 => 7857917,
    234 => 5903370,
    235 => 7173032,
    236 => 3699596,
    237 => 7329447,
    238 => 1341330,
    239 => 4834730,
    240 => 2680103,
    241 => 5187039,
    242 => 126922,
    243 => 4603424,
    244 => 7841118,
    245 => 1595974,
    246 => 7063561,
    247 => 4546524,
    248 => 280005,
    249 => 4784579,
    250 => 6949987,
    251 => 6581310,
    252 => 5582638,
    253 => 6417775,
    254 => 3839961,
    255 => 1976782
  );
-- 256 => 8380416
--   257 => 8378664,
--   258 => 5307408,
--   259 => 1623354,
--   260 => 4778199,
--   261 => 4146264,
--   262 => 2579253,
--   263 => 4385746,
--   264 => 3370349,
--   265 => 27812,
--   266 => 6852351,
--   267 => 3033742,
--   268 => 4965348,
--   269 => 5382198,
--   270 => 7023969,
--   271 => 2185084,
--   272 => 601683,
--   273 => 7198174,
--   274 => 5871437,
--   275 => 1476985,
--   276 => 7986269,
--   277 => 4633167,
--   278 => 1317678,
--   279 => 5274859,
--   280 => 3227876,
--   281 => 1685153,
--   282 => 4166425,
--   283 => 4399818,
--   284 => 2897314,
--   285 => 458740,
--   286 => 8031605,
--   287 => 303005,
--   288 => 3201494,
--   289 => 5720009,
--   290 => 4197045,
--   291 => 7794176,
--   292 => 3110818,
--   293 => 5992904,
--   294 => 4898211,
--   295 => 5016875,
--   296 => 3524442,
--   297 => 1979497,
--   298 => 565603,
--   299 => 2612853,
--   300 => 4623627,
--   301 => 1354892,
--   302 => 3467665,
--   303 => 3014420,
--   304 => 4615550,
--   305 => 3956745,
--   306 => 5569126,
--   307 => 7872490,
--   308 => 6308588,
--   309 => 5184741,
--   310 => 4478945,
--   311 => 7520273,
--   312 => 642628,
--   313 => 3551006,
--   314 => 6644104,
--   315 => 6715099,
--   316 => 5463079,
--   317 => 6341273,
--   318 => 3818627,
--   319 => 6480365,
--   320 => 4614810,
--   321 => 2659525,
--   322 => 2635473,
--   323 => 2374402,
--   324 => 5639874,
--   325 => 6187479,
--   326 => 2391089,
--   327 => 1370517,
--   328 => 5717039,
--   329 => 7371052,
--   330 => 7231559,
--   331 => 5732423,
--   332 => 817536,
--   333 => 89301,
--   334 => 5697147,
--   335 => 6022044,
--   336 => 5698129,
--   337 => 7743490,
--   338 => 6442847,
--   339 => 5889092,
--   340 => 7284949,
--   341 => 7140506,
--   342 => 5344437,
--   343 => 7872272,
--   344 => 5926434,
--   345 => 5702139,
--   346 => 6392603,
--   347 => 1615530,
--   348 => 7823561,
--   349 => 4340221,
--   350 => 7369194,
--   351 => 3974485,
--   352 => 3145678,
--   353 => 59148,
--   354 => 3121440,
--   355 => 7852436,
--   356 => 4675594,
--   357 => 268456,
--   358 => 1300016,
--   359 => 7835041,
--   360 => 7703827,
--   361 => 3956944,
--   362 => 5917973,
--   363 => 7630840,
--   364 => 1716988,
--   365 => 1310261,
--   366 => 653275,
--   367 => 5454363,
--   368 => 7822959,
--   369 => 3284915,
--   370 => 1109516,
--   371 => 724804,
--   372 => 5138445,
--   373 => 7126227,
--   374 => 5454601,
--   375 => 8240173,
--   376 => 5564778,
--   377 => 250446,
--   378 => 3250154,
--   379 => 7216819,
--   380 => 5034454,
--   381 => 818761,
--   382 => 2236726,
--   383 => 7325939,
--   384 => 3572223,
--   385 => 1935420,
--   386 => 7102792,
--   387 => 6275131,
--   388 => 5197539,
--   389 => 1772588,
--   390 => 6592474,
--   391 => 11879,
--   392 => 4063053,
--   393 => 7557876,
--   394 => 7897768,
--   395 => 338420,
--   396 => 6621070,
--   397 => 8238582,
--   398 => 2775755,
--   399 => 5256655,
--   400 => 4837932,
--   401 => 8293209,
--   402 => 6352299,
--   403 => 6386371,
--   404 => 7451668,
--   405 => 6084318,
--   406 => 5919030,
--   407 => 1103344,
--   408 => 6666122,
--   409 => 3410568,
--   410 => 3488383,
--   411 => 5811406,
--   412 => 5188063,
--   413 => 1921994,
--   414 => 327848,
--   415 => 4849188,
--   416 => 2883726,
--   417 => 1780227,
--   418 => 3222807,
--   419 => 1179613,
--   420 => 6279007,
--   421 => 3611750,
--   422 => 4182915,
--   423 => 8165537,
--   424 => 434125,
--   425 => 6783595,
--   426 => 8210729,
--   427 => 4231948,
--   428 => 1935799,
--   429 => 7767179,
--   430 => 6067579,
--   431 => 1716814,
--   432 => 1005239,
--   433 => 2296397,
--   434 => 2983781,
--   435 => 1187885,
--   436 => 4018989,
--   437 => 5737437,
--   438 => 1226661,
--   439 => 4949981,
--   440 => 3585098,
--   441 => 7744461,
--   442 => 8145010,
--   443 => 6352379,
--   444 => 6526611,
--   445 => 1879878,
--   446 => 1922253,
--   447 => 781875,
--   448 => 4618904,
--   449 => 1455890,
--   450 => 4528402,
--   451 => 2033807,
--   452 => 3586446,
--   453 => 1727088,
--   454 => 2254727,
--   455 => 5360024,
--   456 => 1674615,
--   457 => 2454145,
--   458 => 2962264,
--   459 => 5370669,
--   460 => 3574466,
--   461 => 5867399,
--   462 => 2778788,
--   463 => 2193087,
--   464 => 6250525,
--   465 => 3965306,
--   466 => 3815725,
--   467 => 1393159,
--   468 => 3506380,
--   469 => 3838479,
--   470 => 7759253,
--   471 => 553718,
--   472 => 6919699,
--   473 => 3768948,
--   474 => 3197248,
--   475 => 6657188,
--   476 => 4510100,
--   477 => 3472069,
--   478 => 2354215,
--   479 => 3773731,
--   480 => 3201430,
--   481 => 5607817,
--   482 => 274060,
--   483 => 2743411,
--   484 => 7220542,
--   485 => 3180456,
--   486 => 2362063,
--   487 => 770441,
--   488 => 1335936,
--   489 => 3759465,
--   490 => 3334383,
--   491 => 4022750,
--   492 => 3950053,
--   493 => 2218467,
--   494 => 459163,
--   495 => 392707,
--   496 => 1221177,
--   497 => 3716946,
--   498 => 4222329,
--   499 => 1834526,
--   500 => 6224367,
--   501 => 12417,
--   502 => 5006167,
--   503 => 1514152,
--   504 => 6096684,
--   505 => 2455377,
--   506 => 5121960,
--   507 => 3369273,
--   508 => 6522001,
--   509 => 2178965,
--   510 => 6635910,
--   511 => 731434
-- );

end package zeta_lut;
