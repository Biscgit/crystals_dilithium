library work;
  use work.globals.all;

package zeta_lut is

  type zeta_array_t is array (0 to n - 1) of modq_t;

  -- constant zetas : zeta_array_t :=
  -- (
  --   0 => 1,
  --   1 => 42,
  --   2 => 69,
  --   3 => 73,
  --   4 => 15,
  --   5 => 65,
  --   6 => 18,
  --   7 => 78
  -- );

  constant zetas : zeta_array_t :=
  (
    0   => 0,
    1   => 25847,
    2   => 5771523,
    3   => 7861508,
    4   => 237124,
    5   => 7602457,
    6   => 7504169,
    7   => 466468,
    8   => 1826347,
    9   => 2353451,
    10  => 8021166,
    11  => 6288512,
    12  => 3119733,
    13  => 5495562,
    14  => 3111497,
    15  => 2680103,
    16  => 2725464,
    17  => 1024112,
    18  => 7300517,
    19  => 3585928,
    20  => 7830929,
    21  => 7260833,
    22  => 2619752,
    23  => 6271868,
    24  => 6262231,
    25  => 4520680,
    26  => 6980856,
    27  => 5102745,
    28  => 1757237,
    29  => 8360995,
    30  => 4010497,
    31  => 280005,
    32  => 2706023,
    33  => 95776,
    34  => 3077325,
    35  => 3530437,
    36  => 6718724,
    37  => 4788269,
    38  => 5842901,
    39  => 3915439,
    40  => 4519302,
    41  => 5336701,
    42  => 3574422,
    43  => 5512770,
    44  => 3539968,
    45  => 8079950,
    46  => 2348700,
    47  => 7841118,
    48  => 6681150,
    49  => 6736599,
    50  => 3505694,
    51  => 4558682,
    52  => 3507263,
    53  => 6239768,
    54  => 6779997,
    55  => 3699596,
    56  => 811944,
    57  => 531354,
    58  => 954230,
    59  => 3881043,
    60  => 3900724,
    61  => 5823537,
    62  => 2071892,
    63  => 5582638,
    64  => 4450022,
    65  => 6851714,
    66  => 4702672,
    67  => 5339162,
    68  => 6927966,
    69  => 3475950,
    70  => 2176455,
    71  => 6795196,
    72  => 7122806,
    73  => 1939314,
    74  => 4296819,
    75  => 7380215,
    76  => 5190273,
    77  => 5223087,
    78  => 4747489,
    79  => 126922,
    80  => 3412210,
    81  => 7396998,
    82  => 2147896,
    83  => 2715295,
    84  => 5412772,
    85  => 4686924,
    86  => 7969390,
    87  => 5903370,
    88  => 7709315,
    89  => 7151892,
    90  => 8357436,
    91  => 7072248,
    92  => 7998430,
    93  => 1349076,
    94  => 1852771,
    95  => 6949987,
    96  => 5037034,
    97  => 264944,
    98  => 508951,
    99  => 3097992,
    100 => 44288,
    101 => 7280319,
    102 => 904516,
    103 => 3958618,
    104 => 4656075,
    105 => 8371839,
    106 => 1653064,
    107 => 5130689,
    108 => 2389356,
    109 => 8169440,
    110 => 759969,
    111 => 7063561,
    112 => 189548,
    113 => 4827145,
    114 => 3159746,
    115 => 6529015,
    116 => 5971092,
    117 => 8202977,
    118 => 1315589,
    119 => 1341330,
    120 => 1285669,
    121 => 6795489,
    122 => 7567685,
    123 => 6940675,
    124 => 5361315,
    125 => 4499357,
    126 => 4751448,
    127 => 3839961,
    128 => 2091667,
    129 => 3407706,
    130 => 2316500,
    131 => 3817976,
    132 => 5037939,
    133 => 2244091,
    134 => 5933984,
    135 => 4817955,
    136 => 266997,
    137 => 2434439,
    138 => 7144689,
    139 => 3513181,
    140 => 4860065,
    141 => 4621053,
    142 => 7183191,
    143 => 5187039,
    144 => 900702,
    145 => 1859098,
    146 => 909542,
    147 => 819034,
    148 => 495491,
    149 => 6767243,
    150 => 8337157,
    151 => 7857917,
    152 => 7725090,
    153 => 5257975,
    154 => 2031748,
    155 => 3207046,
    156 => 4823422,
    157 => 7855319,
    158 => 7611795,
    159 => 4784579,
    160 => 342297,
    161 => 286988,
    162 => 5942594,
    163 => 4108315,
    164 => 3437287,
    165 => 5038140,
    166 => 1735879,
    167 => 203044,
    168 => 2842341,
    169 => 2691481,
    170 => 5790267,
    171 => 1265009,
    172 => 4055324,
    173 => 1247620,
    174 => 2486353,
    175 => 1595974,
    176 => 4613401,
    177 => 1250494,
    178 => 2635921,
    179 => 4832145,
    180 => 5386378,
    181 => 1869119,
    182 => 1903435,
    183 => 7329447,
    184 => 7047359,
    185 => 1237275,
    186 => 5062207,
    187 => 6950192,
    188 => 7929317,
    189 => 1312455,
    190 => 3306115,
    191 => 6417775,
    192 => 7100756,
    193 => 1917081,
    194 => 5834105,
    195 => 7005614,
    196 => 1500165,
    197 => 777191,
    198 => 2235880,
    199 => 3406031,
    200 => 7838005,
    201 => 5548557,
    202 => 6709241,
    203 => 6533464,
    204 => 5796124,
    205 => 4656147,
    206 => 594136,
    207 => 4603424,
    208 => 6366809,
    209 => 2432395,
    210 => 2454455,
    211 => 8215696,
    212 => 1957272,
    213 => 3369112,
    214 => 185531,
    215 => 7173032,
    216 => 5196991,
    217 => 162844,
    218 => 1616392,
    219 => 3014001,
    220 => 810149,
    221 => 1652634,
    222 => 4686184,
    223 => 6581310,
    224 => 5341501,
    225 => 3523897,
    226 => 3866901,
    227 => 269760,
    228 => 2213111,
    229 => 7404533,
    230 => 1717735,
    231 => 472078,
    232 => 7953734,
    233 => 1723600,
    234 => 6577327,
    235 => 1910376,
    236 => 6712985,
    237 => 7276084,
    238 => 8119771,
    239 => 4546524,
    240 => 5441381,
    241 => 6144432,
    242 => 7959518,
    243 => 6094090,
    244 => 183443,
    245 => 7403526,
    246 => 1612842,
    247 => 4834730,
    248 => 7826001,
    249 => 3919660,
    250 => 8332111,
    251 => 7018208,
    252 => 3937738,
    253 => 1400424,
    254 => 7534263,
    255 => 1976782
  );
-- 256 => 8380416
--   257 => 8378664,
--   258 => 5307408,
--   259 => 1623354,
--   260 => 4778199,
--   261 => 4146264,
--   262 => 2579253,
--   263 => 4385746,
--   264 => 3370349,
--   265 => 27812,
--   266 => 6852351,
--   267 => 3033742,
--   268 => 4965348,
--   269 => 5382198,
--   270 => 7023969,
--   271 => 2185084,
--   272 => 601683,
--   273 => 7198174,
--   274 => 5871437,
--   275 => 1476985,
--   276 => 7986269,
--   277 => 4633167,
--   278 => 1317678,
--   279 => 5274859,
--   280 => 3227876,
--   281 => 1685153,
--   282 => 4166425,
--   283 => 4399818,
--   284 => 2897314,
--   285 => 458740,
--   286 => 8031605,
--   287 => 303005,
--   288 => 3201494,
--   289 => 5720009,
--   290 => 4197045,
--   291 => 7794176,
--   292 => 3110818,
--   293 => 5992904,
--   294 => 4898211,
--   295 => 5016875,
--   296 => 3524442,
--   297 => 1979497,
--   298 => 565603,
--   299 => 2612853,
--   300 => 4623627,
--   301 => 1354892,
--   302 => 3467665,
--   303 => 3014420,
--   304 => 4615550,
--   305 => 3956745,
--   306 => 5569126,
--   307 => 7872490,
--   308 => 6308588,
--   309 => 5184741,
--   310 => 4478945,
--   311 => 7520273,
--   312 => 642628,
--   313 => 3551006,
--   314 => 6644104,
--   315 => 6715099,
--   316 => 5463079,
--   317 => 6341273,
--   318 => 3818627,
--   319 => 6480365,
--   320 => 4614810,
--   321 => 2659525,
--   322 => 2635473,
--   323 => 2374402,
--   324 => 5639874,
--   325 => 6187479,
--   326 => 2391089,
--   327 => 1370517,
--   328 => 5717039,
--   329 => 7371052,
--   330 => 7231559,
--   331 => 5732423,
--   332 => 817536,
--   333 => 89301,
--   334 => 5697147,
--   335 => 6022044,
--   336 => 5698129,
--   337 => 7743490,
--   338 => 6442847,
--   339 => 5889092,
--   340 => 7284949,
--   341 => 7140506,
--   342 => 5344437,
--   343 => 7872272,
--   344 => 5926434,
--   345 => 5702139,
--   346 => 6392603,
--   347 => 1615530,
--   348 => 7823561,
--   349 => 4340221,
--   350 => 7369194,
--   351 => 3974485,
--   352 => 3145678,
--   353 => 59148,
--   354 => 3121440,
--   355 => 7852436,
--   356 => 4675594,
--   357 => 268456,
--   358 => 1300016,
--   359 => 7835041,
--   360 => 7703827,
--   361 => 3956944,
--   362 => 5917973,
--   363 => 7630840,
--   364 => 1716988,
--   365 => 1310261,
--   366 => 653275,
--   367 => 5454363,
--   368 => 7822959,
--   369 => 3284915,
--   370 => 1109516,
--   371 => 724804,
--   372 => 5138445,
--   373 => 7126227,
--   374 => 5454601,
--   375 => 8240173,
--   376 => 5564778,
--   377 => 250446,
--   378 => 3250154,
--   379 => 7216819,
--   380 => 5034454,
--   381 => 818761,
--   382 => 2236726,
--   383 => 7325939,
--   384 => 3572223,
--   385 => 1935420,
--   386 => 7102792,
--   387 => 6275131,
--   388 => 5197539,
--   389 => 1772588,
--   390 => 6592474,
--   391 => 11879,
--   392 => 4063053,
--   393 => 7557876,
--   394 => 7897768,
--   395 => 338420,
--   396 => 6621070,
--   397 => 8238582,
--   398 => 2775755,
--   399 => 5256655,
--   400 => 4837932,
--   401 => 8293209,
--   402 => 6352299,
--   403 => 6386371,
--   404 => 7451668,
--   405 => 6084318,
--   406 => 5919030,
--   407 => 1103344,
--   408 => 6666122,
--   409 => 3410568,
--   410 => 3488383,
--   411 => 5811406,
--   412 => 5188063,
--   413 => 1921994,
--   414 => 327848,
--   415 => 4849188,
--   416 => 2883726,
--   417 => 1780227,
--   418 => 3222807,
--   419 => 1179613,
--   420 => 6279007,
--   421 => 3611750,
--   422 => 4182915,
--   423 => 8165537,
--   424 => 434125,
--   425 => 6783595,
--   426 => 8210729,
--   427 => 4231948,
--   428 => 1935799,
--   429 => 7767179,
--   430 => 6067579,
--   431 => 1716814,
--   432 => 1005239,
--   433 => 2296397,
--   434 => 2983781,
--   435 => 1187885,
--   436 => 4018989,
--   437 => 5737437,
--   438 => 1226661,
--   439 => 4949981,
--   440 => 3585098,
--   441 => 7744461,
--   442 => 8145010,
--   443 => 6352379,
--   444 => 6526611,
--   445 => 1879878,
--   446 => 1922253,
--   447 => 781875,
--   448 => 4618904,
--   449 => 1455890,
--   450 => 4528402,
--   451 => 2033807,
--   452 => 3586446,
--   453 => 1727088,
--   454 => 2254727,
--   455 => 5360024,
--   456 => 1674615,
--   457 => 2454145,
--   458 => 2962264,
--   459 => 5370669,
--   460 => 3574466,
--   461 => 5867399,
--   462 => 2778788,
--   463 => 2193087,
--   464 => 6250525,
--   465 => 3965306,
--   466 => 3815725,
--   467 => 1393159,
--   468 => 3506380,
--   469 => 3838479,
--   470 => 7759253,
--   471 => 553718,
--   472 => 6919699,
--   473 => 3768948,
--   474 => 3197248,
--   475 => 6657188,
--   476 => 4510100,
--   477 => 3472069,
--   478 => 2354215,
--   479 => 3773731,
--   480 => 3201430,
--   481 => 5607817,
--   482 => 274060,
--   483 => 2743411,
--   484 => 7220542,
--   485 => 3180456,
--   486 => 2362063,
--   487 => 770441,
--   488 => 1335936,
--   489 => 3759465,
--   490 => 3334383,
--   491 => 4022750,
--   492 => 3950053,
--   493 => 2218467,
--   494 => 459163,
--   495 => 392707,
--   496 => 1221177,
--   497 => 3716946,
--   498 => 4222329,
--   499 => 1834526,
--   500 => 6224367,
--   501 => 12417,
--   502 => 5006167,
--   503 => 1514152,
--   504 => 6096684,
--   505 => 2455377,
--   506 => 5121960,
--   507 => 3369273,
--   508 => 6522001,
--   509 => 2178965,
--   510 => 6635910,
--   511 => 731434
-- );

end package zeta_lut;
