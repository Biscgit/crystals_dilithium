library work;
  use work.globals.all;

package zeta_lut is

  type zeta_array_t is array (0 to n - 1) of modq_t;

  constant zetas : zeta_array_t :=
  (
    0   => 1,
    1   => 1753,
    2   => 3073009,
    3   => 6757063,
    4   => 3602218,
    5   => 4234153,
    6   => 5801164,
    7   => 3994671,
    8   => 5010068,
    9   => 8352605,
    10  => 1528066,
    11  => 5346675,
    12  => 3415069,
    13  => 2998219,
    14  => 1356448,
    15  => 6195333,
    16  => 7778734,
    17  => 1182243,
    18  => 2508980,
    19  => 6903432,
    20  => 394148,
    21  => 3747250,
    22  => 7062739,
    23  => 3105558,
    24  => 5152541,
    25  => 6695264,
    26  => 4213992,
    27  => 3980599,
    28  => 5483103,
    29  => 7921677,
    30  => 348812,
    31  => 8077412,
    32  => 5178923,
    33  => 2660408,
    34  => 4183372,
    35  => 586241,
    36  => 5269599,
    37  => 2387513,
    38  => 3482206,
    39  => 3363542,
    40  => 4855975,
    41  => 6400920,
    42  => 7814814,
    43  => 5767564,
    44  => 3756790,
    45  => 7025525,
    46  => 4912752,
    47  => 5365997,
    48  => 3764867,
    49  => 4423672,
    50  => 2811291,
    51  => 507927,
    52  => 2071829,
    53  => 3195676,
    54  => 3901472,
    55  => 860144,
    56  => 7737789,
    57  => 4829411,
    58  => 1736313,
    59  => 1665318,
    60  => 2917338,
    61  => 2039144,
    62  => 4561790,
    63  => 1900052,
    64  => 3765607,
    65  => 5720892,
    66  => 5744944,
    67  => 6006015,
    68  => 2740543,
    69  => 2192938,
    70  => 5989328,
    71  => 7009900,
    72  => 2663378,
    73  => 1009365,
    74  => 1148858,
    75  => 2647994,
    76  => 7562881,
    77  => 8291116,
    78  => 2683270,
    79  => 2358373,
    80  => 2682288,
    81  => 636927,
    82  => 1937570,
    83  => 2491325,
    84  => 1095468,
    85  => 1239911,
    86  => 3035980,
    87  => 508145,
    88  => 2453983,
    89  => 2678278,
    90  => 1987814,
    91  => 6764887,
    92  => 556856,
    93  => 4040196,
    94  => 1011223,
    95  => 4405932,
    96  => 5234739,
    97  => 8321269,
    98  => 5258977,
    99  => 527981,
    100 => 3704823,
    101 => 8111961,
    102 => 7080401,
    103 => 545376,
    104 => 676590,
    105 => 4423473,
    106 => 2462444,
    107 => 749577,
    108 => 6663429,
    109 => 7070156,
    110 => 7727142,
    111 => 2926054,
    112 => 557458,
    113 => 5095502,
    114 => 7270901,
    115 => 7655613,
    116 => 3241972,
    117 => 1254190,
    118 => 2925816,
    119 => 140244,
    120 => 2815639,
    121 => 8129971,
    122 => 5130263,
    123 => 1163598,
    124 => 3345963,
    125 => 7561656,
    126 => 6143691,
    127 => 1054478,
    128 => 4808194,
    129 => 6444997,
    130 => 1277625,
    131 => 2105286,
    132 => 3182878,
    133 => 6607829,
    134 => 1787943,
    135 => 8368538,
    136 => 4317364,
    137 => 822541,
    138 => 482649,
    139 => 8041997,
    140 => 1759347,
    141 => 141835,
    142 => 5604662,
    143 => 3123762,
    144 => 3542485,
    145 => 87208,
    146 => 2028118,
    147 => 1994046,
    148 => 928749,
    149 => 2296099,
    150 => 2461387,
    151 => 7277073,
    152 => 1714295,
    153 => 4969849,
    154 => 4892034,
    155 => 2569011,
    156 => 3192354,
    157 => 6458423,
    158 => 8052569,
    159 => 3531229,
    160 => 5496691,
    161 => 6600190,
    162 => 5157610,
    163 => 7200804,
    164 => 2101410,
    165 => 4768667,
    166 => 4197502,
    167 => 214880,
    168 => 7946292,
    169 => 1596822,
    170 => 169688,
    171 => 4148469,
    172 => 6444618,
    173 => 613238,
    174 => 2312838,
    175 => 6663603,
    176 => 7375178,
    177 => 6084020,
    178 => 5396636,
    179 => 7192532,
    180 => 4361428,
    181 => 2642980,
    182 => 7153756,
    183 => 3430436,
    184 => 4795319,
    185 => 635956,
    186 => 235407,
    187 => 2028038,
    188 => 1853806,
    189 => 6500539,
    190 => 6458164,
    191 => 7598542,
    192 => 3761513,
    193 => 6924527,
    194 => 3852015,
    195 => 6346610,
    196 => 4793971,
    197 => 6653329,
    198 => 6125690,
    199 => 3020393,
    200 => 6705802,
    201 => 5926272,
    202 => 5418153,
    203 => 3009748,
    204 => 4805951,
    205 => 2513018,
    206 => 5601629,
    207 => 6187330,
    208 => 2129892,
    209 => 4415111,
    210 => 4564692,
    211 => 6987258,
    212 => 4874037,
    213 => 4541938,
    214 => 621164,
    215 => 7826699,
    216 => 1460718,
    217 => 4611469,
    218 => 5183169,
    219 => 1723229,
    220 => 3870317,
    221 => 4908348,
    222 => 6026202,
    223 => 4606686,
    224 => 5178987,
    225 => 2772600,
    226 => 8106357,
    227 => 5637006,
    228 => 1159875,
    229 => 5199961,
    230 => 6018354,
    231 => 7609976,
    232 => 7044481,
    233 => 4620952,
    234 => 5046034,
    235 => 4357667,
    236 => 4430364,
    237 => 6161950,
    238 => 7921254,
    239 => 7987710,
    240 => 7159240,
    241 => 4663471,
    242 => 4158088,
    243 => 6545891,
    244 => 2156050,
    245 => 8368000,
    246 => 3374250,
    247 => 6866265,
    248 => 2283733,
    249 => 5925040,
    250 => 3258457,
    251 => 5011144,
    252 => 1858416,
    253 => 6201452,
    254 => 1744507,
    255 => 7648983
  );
-- 256 => 8380416
--   257 => 8378664,
--   258 => 5307408,
--   259 => 1623354,
--   260 => 4778199,
--   261 => 4146264,
--   262 => 2579253,
--   263 => 4385746,
--   264 => 3370349,
--   265 => 27812,
--   266 => 6852351,
--   267 => 3033742,
--   268 => 4965348,
--   269 => 5382198,
--   270 => 7023969,
--   271 => 2185084,
--   272 => 601683,
--   273 => 7198174,
--   274 => 5871437,
--   275 => 1476985,
--   276 => 7986269,
--   277 => 4633167,
--   278 => 1317678,
--   279 => 5274859,
--   280 => 3227876,
--   281 => 1685153,
--   282 => 4166425,
--   283 => 4399818,
--   284 => 2897314,
--   285 => 458740,
--   286 => 8031605,
--   287 => 303005,
--   288 => 3201494,
--   289 => 5720009,
--   290 => 4197045,
--   291 => 7794176,
--   292 => 3110818,
--   293 => 5992904,
--   294 => 4898211,
--   295 => 5016875,
--   296 => 3524442,
--   297 => 1979497,
--   298 => 565603,
--   299 => 2612853,
--   300 => 4623627,
--   301 => 1354892,
--   302 => 3467665,
--   303 => 3014420,
--   304 => 4615550,
--   305 => 3956745,
--   306 => 5569126,
--   307 => 7872490,
--   308 => 6308588,
--   309 => 5184741,
--   310 => 4478945,
--   311 => 7520273,
--   312 => 642628,
--   313 => 3551006,
--   314 => 6644104,
--   315 => 6715099,
--   316 => 5463079,
--   317 => 6341273,
--   318 => 3818627,
--   319 => 6480365,
--   320 => 4614810,
--   321 => 2659525,
--   322 => 2635473,
--   323 => 2374402,
--   324 => 5639874,
--   325 => 6187479,
--   326 => 2391089,
--   327 => 1370517,
--   328 => 5717039,
--   329 => 7371052,
--   330 => 7231559,
--   331 => 5732423,
--   332 => 817536,
--   333 => 89301,
--   334 => 5697147,
--   335 => 6022044,
--   336 => 5698129,
--   337 => 7743490,
--   338 => 6442847,
--   339 => 5889092,
--   340 => 7284949,
--   341 => 7140506,
--   342 => 5344437,
--   343 => 7872272,
--   344 => 5926434,
--   345 => 5702139,
--   346 => 6392603,
--   347 => 1615530,
--   348 => 7823561,
--   349 => 4340221,
--   350 => 7369194,
--   351 => 3974485,
--   352 => 3145678,
--   353 => 59148,
--   354 => 3121440,
--   355 => 7852436,
--   356 => 4675594,
--   357 => 268456,
--   358 => 1300016,
--   359 => 7835041,
--   360 => 7703827,
--   361 => 3956944,
--   362 => 5917973,
--   363 => 7630840,
--   364 => 1716988,
--   365 => 1310261,
--   366 => 653275,
--   367 => 5454363,
--   368 => 7822959,
--   369 => 3284915,
--   370 => 1109516,
--   371 => 724804,
--   372 => 5138445,
--   373 => 7126227,
--   374 => 5454601,
--   375 => 8240173,
--   376 => 5564778,
--   377 => 250446,
--   378 => 3250154,
--   379 => 7216819,
--   380 => 5034454,
--   381 => 818761,
--   382 => 2236726,
--   383 => 7325939,
--   384 => 3572223,
--   385 => 1935420,
--   386 => 7102792,
--   387 => 6275131,
--   388 => 5197539,
--   389 => 1772588,
--   390 => 6592474,
--   391 => 11879,
--   392 => 4063053,
--   393 => 7557876,
--   394 => 7897768,
--   395 => 338420,
--   396 => 6621070,
--   397 => 8238582,
--   398 => 2775755,
--   399 => 5256655,
--   400 => 4837932,
--   401 => 8293209,
--   402 => 6352299,
--   403 => 6386371,
--   404 => 7451668,
--   405 => 6084318,
--   406 => 5919030,
--   407 => 1103344,
--   408 => 6666122,
--   409 => 3410568,
--   410 => 3488383,
--   411 => 5811406,
--   412 => 5188063,
--   413 => 1921994,
--   414 => 327848,
--   415 => 4849188,
--   416 => 2883726,
--   417 => 1780227,
--   418 => 3222807,
--   419 => 1179613,
--   420 => 6279007,
--   421 => 3611750,
--   422 => 4182915,
--   423 => 8165537,
--   424 => 434125,
--   425 => 6783595,
--   426 => 8210729,
--   427 => 4231948,
--   428 => 1935799,
--   429 => 7767179,
--   430 => 6067579,
--   431 => 1716814,
--   432 => 1005239,
--   433 => 2296397,
--   434 => 2983781,
--   435 => 1187885,
--   436 => 4018989,
--   437 => 5737437,
--   438 => 1226661,
--   439 => 4949981,
--   440 => 3585098,
--   441 => 7744461,
--   442 => 8145010,
--   443 => 6352379,
--   444 => 6526611,
--   445 => 1879878,
--   446 => 1922253,
--   447 => 781875,
--   448 => 4618904,
--   449 => 1455890,
--   450 => 4528402,
--   451 => 2033807,
--   452 => 3586446,
--   453 => 1727088,
--   454 => 2254727,
--   455 => 5360024,
--   456 => 1674615,
--   457 => 2454145,
--   458 => 2962264,
--   459 => 5370669,
--   460 => 3574466,
--   461 => 5867399,
--   462 => 2778788,
--   463 => 2193087,
--   464 => 6250525,
--   465 => 3965306,
--   466 => 3815725,
--   467 => 1393159,
--   468 => 3506380,
--   469 => 3838479,
--   470 => 7759253,
--   471 => 553718,
--   472 => 6919699,
--   473 => 3768948,
--   474 => 3197248,
--   475 => 6657188,
--   476 => 4510100,
--   477 => 3472069,
--   478 => 2354215,
--   479 => 3773731,
--   480 => 3201430,
--   481 => 5607817,
--   482 => 274060,
--   483 => 2743411,
--   484 => 7220542,
--   485 => 3180456,
--   486 => 2362063,
--   487 => 770441,
--   488 => 1335936,
--   489 => 3759465,
--   490 => 3334383,
--   491 => 4022750,
--   492 => 3950053,
--   493 => 2218467,
--   494 => 459163,
--   495 => 392707,
--   496 => 1221177,
--   497 => 3716946,
--   498 => 4222329,
--   499 => 1834526,
--   500 => 6224367,
--   501 => 12417,
--   502 => 5006167,
--   503 => 1514152,
--   504 => 6096684,
--   505 => 2455377,
--   506 => 5121960,
--   507 => 3369273,
--   508 => 6522001,
--   509 => 2178965,
--   510 => 6635910,
--   511 => 731434
-- );

end package zeta_lut;
