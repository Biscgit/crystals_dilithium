library work;
  use work.globals.all;

package ntt_results is

  type result_array is array (0 to n - 1) of integer;

  type values_array is array (0 to n - 1) of modq_t;

  -- constant values  : values_array := (99, 52, 0, 7, 0, 29, 33, 100);
  -- constant results : result_array := (78, 65, 59, 81, 59, 60, 62, 102);

  constant values : values_array :=
  (
    7038168,
    4193173,
    7085032,
    4158962,
    6012315,
    4013021,
    6115917,
    5928675,
    7075316,
    3937349,
    880280,
    8176627,
    893789,
    6576444,
    6575676,
    4062841,
    3710971,
    5149808,
    1065575,
    5918588,
    4364641,
    689952,
    1916869,
    6961268,
    6476142,
    2322755,
    4863002,
    2774535,
    7422378,
    7301770,
    353514,
    5527476,
    7684287,
    2024372,
    5745435,
    5408524,
    5567492,
    7461918,
    6440578,
    6998354,
    1401800,
    5802268,
    1147043,
    3544123,
    8177658,
    8098622,
    7184480,
    5798167,
    3499537,
    3180042,
    7760119,
    1834143,
    6779626,
    2561220,
    4680899,
    4807684,
    6401056,
    5826255,
    4224689,
    2220705,
    1041151,
    4284304,
    585246,
    920439,
    5894892,
    7349867,
    2648125,
    6105354,
    4970683,
    7221751,
    5794606,
    3179877,
    1696030,
    6389119,
    170417,
    1405103,
    8173756,
    6001883,
    4133800,
    99722,
    710143,
    6949105,
    392949,
    3087718,
    3920539,
    4372622,
    2660684,
    5373427,
    3958297,
    1809743,
    492225,
    2669069,
    1597949,
    7221775,
    3138003,
    1658198,
    5335393,
    5602406,
    3591883,
    543948,
    1568440,
    8928,
    7213845,
    958249,
    1477166,
    7964723,
    4062701,
    1660721,
    3168983,
    6485241,
    1113713,
    7601804,
    4496400,
    3317365,
    6654375,
    8233360,
    5734272,
    8135774,
    5156794,
    3743201,
    5642859,
    6454329,
    1721209,
    1992315,
    3026940,
    35819,
    4479738,
    5200117,
    351763,
    7044062,
    8133687,
    3483585,
    8293122,
    736543,
    2167641,
    6593339,
    3107586,
    869296,
    5848665,
    2358419,
    1771330,
    1919698,
    1461310,
    7319493,
    6648718,
    5597648,
    4748346,
    2941919,
    7772750,
    5429605,
    1089691,
    7874488,
    187620,
    1073537,
    5908902,
    6607566,
    7526371,
    7867037,
    86970,
    8313833,
    1358384,
    4803126,
    6372840,
    2556982,
    5471865,
    5117525,
    3937876,
    5734037,
    7340929,
    4157231,
    7566414,
    5242933,
    596379,
    1522116,
    2053884,
    3150974,
    5620481,
    3180543,
    5904515,
    1061465,
    3730078,
    1696005,
    5667430,
    1538876,
    8016479,
    4726440,
    2521765,
    7866845,
    1899363,
    978766,
    2442645,
    3073770,
    7693369,
    6109986,
    232283,
    7927781,
    4928713,
    416761,
    308970,
    875117,
    7968086,
    5416600,
    717735,
    7798544,
    6958184,
    420021,
    3437489,
    853758,
    3145603,
    4129623,
    5900822,
    1521296,
    1742036,
    1946488,
    5605830,
    5153798,
    7819375,
    689567,
    1370564,
    2832023,
    2769630,
    3499712,
    2899141,
    3738747,
    7509596,
    3320067,
    5332485,
    1047449,
    3626703,
    7950452,
    3498218,
    8334557,
    2824960,
    4951468,
    6182818,
    3037921,
    1405326,
    5628031,
    7257637,
    2765458,
    8075481,
    6991205,
    931076,
    5479086,
    8204517,
    6774417,
    4554010,
    2156255,
    7327438,
    3394746,
    418868,
    7287118,
    8343692,
    7657108,
    8349009,
    5574367
  );

  constant results : result_array :=
  (
    3527686,
    1930588,
    3109133,
    5864302,
    5046357,
    7180728,
    3677363,
    7402123,
    5452393,
    3068822,
    4177592,
    3754672,
    6441119,
    834830,
    5593069,
    1346096,
    7433690,
    5248240,
    7381866,
    5971261,
    2848352,
    7529224,
    2276516,
    3969301,
    6655674,
    4238398,
    5688288,
    578381,
    3165083,
    2101219,
    1859125,
    350328,
    1444633,
    7300910,
    825594,
    6641300,
    4108858,
    2293463,
    8138518,
    5193831,
    6105516,
    8002591,
    3579763,
    2793597,
    6321434,
    5400270,
    2649898,
    3691205,
    2584629,
    6544632,
    3227508,
    1259002,
    2295618,
    8102371,
    1360611,
    8073986,
    1865209,
    3686036,
    7018127,
    90248,
    4184999,
    3178362,
    6316209,
    942974,
    7598964,
    715087,
    4306691,
    4000008,
    3941721,
    1634590,
    7963527,
    3320444,
    6674293,
    1141916,
    6067728,
    5018938,
    2639694,
    737792,
    1519410,
    2308218,
    3486301,
    7925840,
    257492,
    1159264,
    3014871,
    8339346,
    6435658,
    8272944,
    2746133,
    4855141,
    6830334,
    358101,
    6965575,
    3249763,
    3852118,
    2963416,
    5103527,
    5083259,
    6246892,
    2527734,
    292616,
    3079781,
    2297553,
    435031,
    1622203,
    208731,
    6995597,
    3110387,
    6129298,
    3534259,
    5385553,
    7385850,
    3809136,
    1280785,
    491589,
    1234377,
    4131310,
    6398603,
    7637128,
    6716713,
    8351908,
    3833405,
    4218043,
    5270090,
    4490416,
    1423582,
    3299068,
    2746643,
    1431861,
    5157381,
    3314567,
    7570866,
    4740801,
    7575541,
    7318172,
    4174501,
    6127722,
    584320,
    4093870,
    1041095,
    352307,
    820593,
    4435463,
    6813754,
    223597,
    1660151,
    1345453,
    7490166,
    1161820,
    8198582,
    3881731,
    6440531,
    7650119,
    1569674,
    6292111,
    432814,
    2351228,
    3023258,
    7437575,
    1195476,
    3735152,
    1483424,
    4480029,
    5156627,
    1057805,
    3022359,
    7248927,
    1355602,
    1804737,
    680166,
    215020,
    1734798,
    3810080,
    8142052,
    7684391,
    820393,
    7490854,
    3634292,
    7457280,
    112414,
    3780885,
    6257111,
    2185076,
    3696558,
    7172198,
    5071839,
    5212423,
    8256215,
    1126156,
    6741083,
    7271950,
    5410663,
    987434,
    680684,
    7655449,
    4178692,
    8222360,
    2038722,
    2199954,
    1146935,
    4442265,
    7197356,
    5108430,
    7688998,
    4752779,
    6964992,
    448449,
    1239143,
    5939096,
    801295,
    1187578,
    6251498,
    7089901,
    5069566,
    3271164,
    4319075,
    6107991,
    7353098,
    3184631,
    4876982,
    255170,
    5011433,
    245355,
    6446093,
    7096027,
    3637946,
    5019147,
    6567199,
    5165127,
    2891287,
    1746549,
    1853072,
    8016272,
    94745,
    8050390,
    6746713,
    2050347,
    863793,
    7467259,
    5434527,
    7126217,
    594550,
    4873370,
    2907134,
    6448770,
    2781075,
    4155076,
    868921,
    995631,
    6152978,
    7846396,
    5934588,
    3419660,
    3415933,
    2593000,
    5525863
  );

end package ntt_results;
