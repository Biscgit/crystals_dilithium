library work;
  use work.globals.all;

package ntt_results is

  type result_array is array (0 to n - 1) of integer;

  type values_array is array (0 to n - 1) of modq_t;

  constant values  : values_array := (99, 52, 0, 7, 0, 29, 33, 100);
  constant results : result_array := (78, 65, 59, 81, 59, 60, 62, 102);

--   constant values : values_array :=
--   (
--     5204207,
--     3889113,
--     6812016,
--     2160869,
--     7641924,
--     6900026,
--     2352012,
--     4919756,
--     5592427,
--     4574255,
--     2033669,
--     4861918,
--     4387486,
--     1127877,
--     5330363,
--     4990563,
--     8291416,
--     5405970,
--     4685707,
--     4311714,
--     7105922,
--     6254811,
--     1257539,
--     1130323,
--     5382954,
--     1283377,
--     3083648,
--     5125843,
--     142388,
--     1546691,
--     1059490,
--     4147902,
--     6119954,
--     1486753,
--     1432834,
--     157027,
--     2722529,
--     2980305,
--     7850180,
--     242830,
--     767456,
--     409707,
--     4889189,
--     3625838,
--     4043404,
--     1705939,
--     8233920,
--     1048147,
--     770380,
--     6679964,
--     6871839,
--     2743704,
--     7274976,
--     3641934,
--     3392294,
--     6488652,
--     2949607,
--     468179,
--     4367368,
--     4715262,
--     4421437,
--     3005143,
--     3967619,
--     982474,
--     4428638,
--     4329653,
--     959570,
--     6007260,
--     8056737,
--     2907741,
--     6850243,
--     446393,
--     7161304,
--     4826340,
--     6327163,
--     7769262,
--     7019287,
--     4666037,
--     2661325,
--     3545364,
--     5522831,
--     3763597,
--     7549150,
--     1805101,
--     3369865,
--     6012623,
--     3230366,
--     7772708,
--     900301,
--     8109643,
--     3539627,
--     6124401,
--     8320059,
--     157533,
--     5273277,
--     1349842,
--     8347996,
--     7696767,
--     3124219,
--     1452430,
--     4126919,
--     7713915,
--     3787057,
--     934543,
--     4636711,
--     916620,
--     4272609,
--     5548821,
--     129508,
--     1882054,
--     2770397,
--     4901514,
--     1709611,
--     605457,
--     4383247,
--     6917574,
--     6799946,
--     1635791,
--     1005873,
--     2374736,
--     6477192,
--     7613984,
--     4712784,
--     4339851,
--     2351150,
--     1833482,
--     306439,
--     6123938,
--     580074,
--     232319,
--     6137619,
--     1811058,
--     5471159,
--     5624568,
--     1242408,
--     972364,
--     4564669,
--     3649647,
--     5249478,
--     4117785,
--     1832797,
--     3913034,
--     3056974,
--     7074006,
--     7338082,
--     8198398,
--     1250144,
--     7033028,
--     892011,
--     6383588,
--     6722645,
--     8071579,
--     4398982,
--     5769656,
--     8034782,
--     4853295,
--     329506,
--     7094037,
--     6629990,
--     3814258,
--     6306447,
--     832717,
--     1436517,
--     3218644,
--     7606694,
--     635192,
--     2847190,
--     207398,
--     6142075,
--     7770030,
--     4190566,
--     2296811,
--     2038267,
--     7682766,
--     5336117,
--     2234254,
--     6409366,
--     7932291,
--     7924866,
--     6355475,
--     6070909,
--     1645687,
--     6657272,
--     6236339,
--     3428304,
--     5757813,
--     7824531,
--     3954450,
--     4385428,
--     4747656,
--     6732377,
--     7855087,
--     4567118,
--     3183387,
--     6811273,
--     2063699,
--     7123619,
--     2519971,
--     1771585,
--     7042975,
--     1042906,
--     4938322,
--     7103735,
--     3393164,
--     2554537,
--     6068816,
--     4381180,
--     7531739,
--     5937445,
--     3628340,
--     3711855,
--     1083202,
--     6524045,
--     1225976,
--     832941,
--     726408,
--     4746057,
--     90229,
--     1725109,
--     4468709,
--     5711664,
--     5858031,
--     6505659,
--     1562067,
--     3494813,
--     1053302,
--     6364852,
--     3436883,
--     2109271,
--     2077737,
--     1069722,
--     667661,
--     931556,
--     5892346,
--     4114175,
--     1078948,
--     7356497,
--     4422717,
--     5443976,
--     6105719,
--     5267639,
--     6560589,
--     5608252,
--     1418728,
--     1829915,
--     794680,
--     3833087,
--     7022285,
--     1725602,
--     8223508,
--     4106720,
--     4465275,
--     1421866,
--     3100798,
--     3906643,
--     2661727
--   );
--
--   constant results : result_array :=
--   (
--     1580717,
--     3208715,
--     - 4732436,
--     2085725,
--     - 2890030,
--     1952753,
--     - 1805438,
--     - 206911,
--     - 6151337,
--     - 2267525,
--     1206187,
--     989810,
--     934374,
--     - 541327,
--     - 2459137,
--     2008675,
--     - 2112143,
--     - 713173,
--     2899539,
--     1786363,
--     - 3294060,
--     - 3592275,
--     5172785,
--     - 313889,
--     4866533,
--     768362,
--     - 2367803,
--     - 2299935,
--     - 1739499,
--     - 34208,
--     - 1091290,
--     - 2481685,
--     - 2684955,
--     1988155,
--     2445999,
--     292220,
--     - 8714056,
--     1942629,
--     - 2534952,
--     1811582,
--     4586767,
--     - 2489045,
--     2312169,
--     3957150,
--     89699,
--     2200588,
--     1722255,
--     - 3096226,
--     3557569,
--     2657848,
--     1848077,
--     - 159826,
--     1087811,
--     678691,
--     3207886,
--     - 4071937,
--     - 2406250,
--     - 734971,
--     - 2993257,
--     4129518,
--     - 5705475,
--     - 1281514,
--     3410267,
--     - 496877,
--     12214381,
--     987447,
--     - 1737484,
--     - 3679598,
--     3116371,
--     2756412,
--     1141562,
--     - 4068692,
--     265445,
--     - 947082,
--     - 6970539,
--     1403022,
--     - 4521379,
--     - 935508,
--     2668994,
--     3411023,
--     3734616,
--     - 2976145,
--     362986,
--     - 1994794,
--     4420015,
--     673130,
--     - 535113,
--     1108358,
--     - 1141891,
--     1762240,
--     188830,
--     - 31651,
--     959353,
--     3195206,
--     4902832,
--     2105012,
--     4873726,
--     - 61440,
--     2716295,
--     3293097,
--     492434,
--     - 3756402,
--     793020,
--     - 3518736,
--     - 2491569,
--     2916109,
--     - 2978229,
--     438508,
--     3039257,
--     - 4042320,
--     - 5381356,
--     1634974,
--     - 10616109,
--     2061910,
--     - 2680220,
--     3431656,
--     339092,
--     422808,
--     1264413,
--     2684895,
--     - 1366933,
--     4176391,
--     - 2155772,
--     131718,
--     - 1130600,
--     - 1267891,
--     422529,
--     136107,
--     - 7940655,
--     546740,
--     - 4893867,
--     - 2132258,
--     - 282208,
--     - 2158930,
--     - 1862940,
--     453118,
--     - 7189984,
--     1004412,
--     - 2750547,
--     - 3130817,
--     - 4094793,
--     - 2875123,
--     - 1540612,
--     - 913724,
--     - 2140286,
--     4046455,
--     - 1853760,
--     3828442,
--     3625224,
--     3718209,
--     693038,
--     - 1424327,
--     - 2139850,
--     - 457067,
--     - 1037487,
--     - 1203038,
--     - 228495,
--     3026743,
--     - 5089927,
--     - 2752728,
--     2751913,
--     - 2531569,
--     368560,
--     1406404,
--     2399163,
--     - 1612023,
--     - 1101387,
--     - 541948,
--     3447425,
--     - 2219041,
--     4413173,
--     205006,
--     6772648,
--     796155,
--     6141341,
--     111603,
--     - 7621833,
--     1841566,
--     3350454,
--     - 1359013,
--     - 8257664,
--     110676,
--     292119,
--     1101359,
--     - 3611572,
--     - 1570118,
--     3640611,
--     - 2362401,
--     - 1724738,
--     3585660,
--     3233173,
--     - 1547735,
--     - 787871,
--     1438771,
--     4067998,
--     2847278,
--     - 509025,
--     - 3964385,
--     - 1085779,
--     3712116,
--     7352880,
--     4053510,
--     2785817,
--     2062577,
--     - 4399186,
--     - 3765660,
--     - 1831674,
--     - 95023,
--     1225942,
--     16030,
--     - 4890473,
--     1993145,
--     1867345,
--     - 3308644,
--     5774808,
--     - 1798969,
--     - 2357907,
--     - 860413,
--     7215080,
--     - 2142384,
--     5461374,
--     - 217880,
--     - 537536,
--     3536332,
--     5911598,
--     - 1829954,
--     642582,
--     1961778,
--     4562454,
--     2416489,
--     926750,
--     2942442,
--     11450259,
--     4059124,
--     - 5137515,
--     - 2908514,
--     1141341,
--     3696519,
--     30833,
--     1227122,
--     - 4761525,
--     - 1861905,
--     - 2475613,
--     3236577,
--     43772,
--     3933149,
--     - 7264071,
--     - 3335729,
--     588657,
--     - 901036,
--     - 25442,
--     1037214,
--     - 1282519,
--     2622412,
--     - 3119293,
--     3644026
--   );
--

end package ntt_results;
